interface adder_if;
    logic       clk;
    logic       rstn;
    logic [4:0] a;
    logic [4:0] b;
    logic [5:0] y;
endinterface