interface dff_if(input bit clk);
    logic rstn;
    logic d;
    logic q;
endinterface